module production (a, b, out0, out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12, out13, out14, out15, out16, out17, out18);
	input[9:0] a;
	input[9:0] b;
	output out0;
	output[1:0] out1;
	output[2:0] out2;
	output[3:0] out3;
	output[4:0] out4;
	output[5:0] out5;
	output[6:0] out6;
	output[7:0] out7;
	output[8:0] out8;
	output[9:0] out9;
	output[8:0] out10;
	output[7:0] out11;
	output[6:0] out12;
	output[5:0] out13;
	output[4:0] out14;
	output[3:0] out15;
	output[2:0] out16;
	output[1:0] out17;
	output out18;
	assign out0 = a[9] & b[9];
	assign out1[0] = a[8] & b[9];
	assign out1[1] = a[9] & b[8];
	assign out2[0] = a[7] & b[9];
	assign out2[1] = a[8] & b[8];
	assign out2[2] = a[9] & b[7];
	assign out3[0] = a[6] & b[9];
	assign out3[1] = a[7] & b[8];
	assign out3[2] = a[8] & b[7];
	assign out3[3] = a[9] & b[6];
	assign out4[0] = a[5] & b[9];
	assign out4[1] = a[6] & b[8];
	assign out4[2] = a[7] & b[7];
	assign out4[3] = a[8] & b[6];
	assign out4[4] = a[9] & b[5];
	assign out5[0] = a[4] & b[9];
	assign out5[1] = a[5] & b[8];
	assign out5[2] = a[6] & b[7];
	assign out5[3] = a[7] & b[6];
	assign out5[4] = a[8] & b[5];
	assign out5[5] = a[9] & b[4];
	assign out6[0] = a[3] & b[9];
	assign out6[1] = a[4] & b[8];
	assign out6[2] = a[5] & b[7];
	assign out6[3] = a[6] & b[6];
	assign out6[4] = a[7] & b[5];
	assign out6[5] = a[8] & b[4];
	assign out6[6] = a[9] & b[3];
	assign out7[0] = a[2] & b[9];
	assign out7[1] = a[3] & b[8];
	assign out7[2] = a[4] & b[7];
	assign out7[3] = a[5] & b[6];
	assign out7[4] = a[6] & b[5];
	assign out7[5] = a[7] & b[4];
	assign out7[6] = a[8] & b[3];
	assign out7[7] = a[9] & b[2];
	assign out8[0] = a[1] & b[9];
	assign out8[1] = a[2] & b[8];
	assign out8[2] = a[3] & b[7];
	assign out8[3] = a[4] & b[6];
	assign out8[4] = a[5] & b[5];
	assign out8[5] = a[6] & b[4];
	assign out8[6] = a[7] & b[3];
	assign out8[7] = a[8] & b[2];
	assign out8[8] = a[9] & b[1];
	assign out9[0] = a[0] & b[9];
	assign out9[1] = a[1] & b[8];
	assign out9[2] = a[2] & b[7];
	assign out9[3] = a[3] & b[6];
	assign out9[4] = a[4] & b[5];
	assign out9[5] = a[5] & b[4];
	assign out9[6] = a[6] & b[3];
	assign out9[7] = a[7] & b[2];
	assign out9[8] = a[8] & b[1];
	assign out9[9] = a[9] & b[0];
	assign out10[0] = a[0] & b[8];
	assign out10[1] = a[1] & b[7];
	assign out10[2] = a[2] & b[6];
	assign out10[3] = a[3] & b[5];
	assign out10[4] = a[4] & b[4];
	assign out10[5] = a[5] & b[3];
	assign out10[6] = a[6] & b[2];
	assign out10[7] = a[7] & b[1];
	assign out10[8] = a[8] & b[0];
	assign out11[0] = a[0] & b[7];
	assign out11[1] = a[1] & b[6];
	assign out11[2] = a[2] & b[5];
	assign out11[3] = a[3] & b[4];
	assign out11[4] = a[4] & b[3];
	assign out11[5] = a[5] & b[2];
	assign out11[6] = a[6] & b[1];
	assign out11[7] = a[7] & b[0];
	assign out12[0] = a[0] & b[6];
	assign out12[1] = a[1] & b[5];
	assign out12[2] = a[2] & b[4];
	assign out12[3] = a[3] & b[3];
	assign out12[4] = a[4] & b[2];
	assign out12[5] = a[5] & b[1];
	assign out12[6] = a[6] & b[0];
	assign out13[0] = a[0] & b[5];
	assign out13[1] = a[1] & b[4];
	assign out13[2] = a[2] & b[3];
	assign out13[3] = a[3] & b[2];
	assign out13[4] = a[4] & b[1];
	assign out13[5] = a[5] & b[0];
	assign out14[0] = a[0] & b[4];
	assign out14[1] = a[1] & b[3];
	assign out14[2] = a[2] & b[2];
	assign out14[3] = a[3] & b[1];
	assign out14[4] = a[4] & b[0];
	assign out15[0] = a[0] & b[3];
	assign out15[1] = a[1] & b[2];
	assign out15[2] = a[2] & b[1];
	assign out15[3] = a[3] & b[0];
	assign out16[0] = a[0] & b[2];
	assign out16[1] = a[1] & b[1];
	assign out16[2] = a[2] & b[0];
	assign out17[0] = a[0] & b[1];
	assign out17[1] = a[1] & b[0];
	assign out18 = a[0] & b[0];
endmodule
