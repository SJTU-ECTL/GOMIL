module Inf2 (a, p, g);
	input a;
	output p;
	output g;
	assign p = a;
	assign g = 0;
endmodule
