module Compress_Tree (a, b, data0_s5, data1_s5, data2_s5, data3_s5, data4_s5, data5_s5, data6_s5, data7_s5, data8_s5, data9_s5, data10_s5, data11_s5, data12_s5, data13_s5, data14_s5, data15_s5, data16_s5, data17_s5, data18_s5);
	input[9:0] a;
	input[9:0] b;
	output[1:0] data0_s5;
	output[1:0] data1_s5;
	output[1:0] data2_s5;
	output[1:0] data3_s5;
	output[1:0] data4_s5;
	output[1:0] data5_s5;
	output[1:0] data6_s5;
	output[1:0] data7_s5;
	output[1:0] data8_s5;
	output[1:0] data9_s5;
	output[1:0] data10_s5;
	output[0:0] data11_s5;
	output[0:0] data12_s5;
	output[1:0] data13_s5;
	output[0:0] data14_s5;
	output[0:0] data15_s5;
	output[0:0] data16_s5;
	output[0:0] data17_s5;
	output[0:0] data18_s5;

	//pre-processing block : production
	wire[0:0] out0;
	wire[1:0] out1;
	wire[2:0] out2;
	wire[3:0] out3;
	wire[4:0] out4;
	wire[5:0] out5;
	wire[6:0] out6;
	wire[7:0] out7;
	wire[8:0] out8;
	wire[9:0] out9;
	wire[8:0] out10;
	wire[7:0] out11;
	wire[6:0] out12;
	wire[5:0] out13;
	wire[4:0] out14;
	wire[3:0] out15;
	wire[2:0] out16;
	wire[1:0] out17;
	wire[0:0] out18;
	production PD0(.a(a),.b(b),.out0(out0),.out1(out1),.out2(out2),.out3(out3),.out4(out4),.out5(out5),.out6(out6),.out7(out7),.out8(out8),.out9(out9),.out10(out10),.out11(out11),.out12(out12),.out13(out13),.out14(out14),.out15(out15),.out16(out16),.out17(out17),.out18(out18));


	//****The 1th stage****
	wire[0:0] data0_s1;
	wire[1:0] data1_s1;
	wire[2:0] data2_s1;
	wire[4:0] data3_s1;
	wire[4:0] data4_s1;
	wire[3:0] data5_s1;
	wire[2:0] data6_s1;
	wire[10:0] data7_s1;
	wire[5:0] data8_s1;
	wire[6:0] data9_s1;
	wire[2:0] data10_s1;
	wire[7:0] data11_s1;
	wire[8:0] data12_s1;
	wire[3:0] data13_s1;
	wire[2:0] data14_s1;
	wire[3:0] data15_s1;
	wire[2:0] data16_s1;
	wire[0:0] data17_s1;
	wire[0:0] data18_s1;
	assign data0_s1[0] = out0[0];
	assign data1_s1[0] = out1[0];
	assign data1_s1[1] = out1[1];
	assign data2_s1[0] = out2[0];
	assign data2_s1[1] = out2[1];
	assign data2_s1[2] = out2[2];
	assign data3_s1[0] = out3[0];
	assign data3_s1[1] = out3[1];
	assign data3_s1[2] = out3[2];
	assign data3_s1[3] = out3[3];
	FA F0(.a(out4[0]),.b(out4[1]),.cin(out4[2]),.sum(data4_s1[0]),.cout(data3_s1[4]));
	assign data4_s1[1] = out4[3];
	assign data4_s1[2] = out4[4];
	FA F1(.a(out5[0]),.b(out5[1]),.cin(out5[2]),.sum(data5_s1[0]),.cout(data4_s1[3]));
	FA F2(.a(out5[3]),.b(out5[4]),.cin(out5[5]),.sum(data5_s1[1]),.cout(data4_s1[4]));
	FA F3(.a(out6[0]),.b(out6[1]),.cin(out6[2]),.sum(data6_s1[0]),.cout(data5_s1[2]));
	FA F4(.a(out6[3]),.b(out6[4]),.cin(out6[5]),.sum(data6_s1[1]),.cout(data5_s1[3]));
	assign data6_s1[2] = out6[6];
	assign data7_s1[0] = out7[0];
	assign data7_s1[1] = out7[1];
	assign data7_s1[2] = out7[2];
	assign data7_s1[3] = out7[3];
	assign data7_s1[4] = out7[4];
	assign data7_s1[5] = out7[5];
	assign data7_s1[6] = out7[6];
	assign data7_s1[7] = out7[7];
	FA F5(.a(out8[0]),.b(out8[1]),.cin(out8[2]),.sum(data8_s1[0]),.cout(data7_s1[8]));
	FA F6(.a(out8[3]),.b(out8[4]),.cin(out8[5]),.sum(data8_s1[1]),.cout(data7_s1[9]));
	FA F7(.a(out8[6]),.b(out8[7]),.cin(out8[8]),.sum(data8_s1[2]),.cout(data7_s1[10]));
	FA F8(.a(out9[0]),.b(out9[1]),.cin(out9[2]),.sum(data9_s1[0]),.cout(data8_s1[3]));
	FA F9(.a(out9[3]),.b(out9[4]),.cin(out9[5]),.sum(data9_s1[1]),.cout(data8_s1[4]));
	FA F10(.a(out9[6]),.b(out9[7]),.cin(out9[8]),.sum(data9_s1[2]),.cout(data8_s1[5]));
	assign data9_s1[3] = out9[9];
	FA F11(.a(out10[0]),.b(out10[1]),.cin(out10[2]),.sum(data10_s1[0]),.cout(data9_s1[4]));
	FA F12(.a(out10[3]),.b(out10[4]),.cin(out10[5]),.sum(data10_s1[1]),.cout(data9_s1[5]));
	FA F13(.a(out10[6]),.b(out10[7]),.cin(out10[8]),.sum(data10_s1[2]),.cout(data9_s1[6]));
	assign data11_s1[0] = out11[0];
	assign data11_s1[1] = out11[1];
	assign data11_s1[2] = out11[2];
	assign data11_s1[3] = out11[3];
	assign data11_s1[4] = out11[4];
	assign data11_s1[5] = out11[5];
	assign data11_s1[6] = out11[6];
	assign data11_s1[7] = out11[7];
	assign data12_s1[0] = out12[0];
	assign data12_s1[1] = out12[1];
	assign data12_s1[2] = out12[2];
	assign data12_s1[3] = out12[3];
	assign data12_s1[4] = out12[4];
	assign data12_s1[5] = out12[5];
	assign data12_s1[6] = out12[6];
	FA F14(.a(out13[0]),.b(out13[1]),.cin(out13[2]),.sum(data13_s1[0]),.cout(data12_s1[7]));
	FA F15(.a(out13[3]),.b(out13[4]),.cin(out13[5]),.sum(data13_s1[1]),.cout(data12_s1[8]));
	FA F16(.a(out14[0]),.b(out14[1]),.cin(out14[2]),.sum(data14_s1[0]),.cout(data13_s1[2]));
	HA H0(.a(out14[3]),.cin(out14[4]),.sum(data14_s1[1]),.cout(data13_s1[3]));
	HA H1(.a(out15[0]),.cin(out15[1]),.sum(data15_s1[0]),.cout(data14_s1[2]));
	assign data15_s1[1] = out15[2];
	assign data15_s1[2] = out15[3];
	HA H2(.a(out16[0]),.cin(out16[1]),.sum(data16_s1[0]),.cout(data15_s1[3]));
	assign data16_s1[1] = out16[2];
	HA H3(.a(out17[0]),.cin(out17[1]),.sum(data17_s1[0]),.cout(data16_s1[2]));
	assign data18_s1[0] = out18[0];

	//****The 2th stage****
	wire[0:0] data0_s2;
	wire[2:0] data1_s2;
	wire[0:0] data2_s2;
	wire[5:0] data3_s2;
	wire[2:0] data4_s2;
	wire[3:0] data5_s2;
	wire[5:0] data6_s2;
	wire[6:0] data7_s2;
	wire[3:0] data8_s2;
	wire[2:0] data9_s2;
	wire[4:0] data10_s2;
	wire[5:0] data11_s2;
	wire[5:0] data12_s2;
	wire[2:0] data13_s2;
	wire[0:0] data14_s2;
	wire[4:0] data15_s2;
	wire[0:0] data16_s2;
	wire[0:0] data17_s2;
	wire[0:0] data18_s2;
	assign data0_s2[0] = data0_s1[0];
	assign data1_s2[0] = data1_s1[0];
	assign data1_s2[1] = data1_s1[1];
	FA F17(.a(data2_s1[0]),.b(data2_s1[1]),.cin(data2_s1[2]),.sum(data2_s2[0]),.cout(data1_s2[2]));
	assign data3_s2[0] = data3_s1[0];
	assign data3_s2[1] = data3_s1[1];
	assign data3_s2[2] = data3_s1[2];
	assign data3_s2[3] = data3_s1[3];
	assign data3_s2[4] = data3_s1[4];
	FA F18(.a(data4_s1[0]),.b(data4_s1[1]),.cin(data4_s1[2]),.sum(data4_s2[0]),.cout(data3_s2[5]));
	assign data4_s2[1] = data4_s1[3];
	assign data4_s2[2] = data4_s1[4];
	assign data5_s2[0] = data5_s1[0];
	assign data5_s2[1] = data5_s1[1];
	assign data5_s2[2] = data5_s1[2];
	assign data5_s2[3] = data5_s1[3];
	assign data6_s2[0] = data6_s1[0];
	assign data6_s2[1] = data6_s1[1];
	assign data6_s2[2] = data6_s1[2];
	FA F19(.a(data7_s1[0]),.b(data7_s1[1]),.cin(data7_s1[2]),.sum(data7_s2[0]),.cout(data6_s2[3]));
	FA F20(.a(data7_s1[3]),.b(data7_s1[4]),.cin(data7_s1[5]),.sum(data7_s2[1]),.cout(data6_s2[4]));
	FA F21(.a(data7_s1[6]),.b(data7_s1[7]),.cin(data7_s1[8]),.sum(data7_s2[2]),.cout(data6_s2[5]));
	assign data7_s2[3] = data7_s1[9];
	assign data7_s2[4] = data7_s1[10];
	FA F22(.a(data8_s1[0]),.b(data8_s1[1]),.cin(data8_s1[2]),.sum(data8_s2[0]),.cout(data7_s2[5]));
	FA F23(.a(data8_s1[3]),.b(data8_s1[4]),.cin(data8_s1[5]),.sum(data8_s2[1]),.cout(data7_s2[6]));
	FA F24(.a(data9_s1[0]),.b(data9_s1[1]),.cin(data9_s1[2]),.sum(data9_s2[0]),.cout(data8_s2[2]));
	FA F25(.a(data9_s1[3]),.b(data9_s1[4]),.cin(data9_s1[5]),.sum(data9_s2[1]),.cout(data8_s2[3]));
	assign data9_s2[2] = data9_s1[6];
	assign data10_s2[0] = data10_s1[0];
	assign data10_s2[1] = data10_s1[1];
	assign data10_s2[2] = data10_s1[2];
	FA F26(.a(data11_s1[0]),.b(data11_s1[1]),.cin(data11_s1[2]),.sum(data11_s2[0]),.cout(data10_s2[3]));
	FA F27(.a(data11_s1[3]),.b(data11_s1[4]),.cin(data11_s1[5]),.sum(data11_s2[1]),.cout(data10_s2[4]));
	assign data11_s2[2] = data11_s1[6];
	assign data11_s2[3] = data11_s1[7];
	FA F28(.a(data12_s1[0]),.b(data12_s1[1]),.cin(data12_s1[2]),.sum(data12_s2[0]),.cout(data11_s2[4]));
	FA F29(.a(data12_s1[3]),.b(data12_s1[4]),.cin(data12_s1[5]),.sum(data12_s2[1]),.cout(data11_s2[5]));
	assign data12_s2[2] = data12_s1[6];
	assign data12_s2[3] = data12_s1[7];
	assign data12_s2[4] = data12_s1[8];
	FA F30(.a(data13_s1[0]),.b(data13_s1[1]),.cin(data13_s1[2]),.sum(data13_s2[0]),.cout(data12_s2[5]));
	assign data13_s2[1] = data13_s1[3];
	FA F31(.a(data14_s1[0]),.b(data14_s1[1]),.cin(data14_s1[2]),.sum(data14_s2[0]),.cout(data13_s2[2]));
	assign data15_s2[0] = data15_s1[0];
	assign data15_s2[1] = data15_s1[1];
	assign data15_s2[2] = data15_s1[2];
	assign data15_s2[3] = data15_s1[3];
	FA F32(.a(data16_s1[0]),.b(data16_s1[1]),.cin(data16_s1[2]),.sum(data16_s2[0]),.cout(data15_s2[4]));
	assign data17_s2[0] = data17_s1[0];
	assign data18_s2[0] = data18_s1[0];

	//****The 3th stage****
	wire[0:0] data0_s3;
	wire[2:0] data1_s3;
	wire[2:0] data2_s3;
	wire[1:0] data3_s3;
	wire[2:0] data4_s3;
	wire[5:0] data5_s3;
	wire[3:0] data6_s3;
	wire[3:0] data7_s3;
	wire[2:0] data8_s3;
	wire[3:0] data9_s3;
	wire[3:0] data10_s3;
	wire[3:0] data11_s3;
	wire[2:0] data12_s3;
	wire[0:0] data13_s3;
	wire[1:0] data14_s3;
	wire[2:0] data15_s3;
	wire[0:0] data16_s3;
	wire[0:0] data17_s3;
	wire[0:0] data18_s3;
	assign data0_s3[0] = data0_s2[0];
	assign data1_s3[0] = data1_s2[0];
	assign data1_s3[1] = data1_s2[1];
	assign data1_s3[2] = data1_s2[2];
	assign data2_s3[0] = data2_s2[0];
	FA F33(.a(data3_s2[0]),.b(data3_s2[1]),.cin(data3_s2[2]),.sum(data3_s3[0]),.cout(data2_s3[1]));
	FA F34(.a(data3_s2[3]),.b(data3_s2[4]),.cin(data3_s2[5]),.sum(data3_s3[1]),.cout(data2_s3[2]));
	assign data4_s3[0] = data4_s2[0];
	assign data4_s3[1] = data4_s2[1];
	assign data4_s3[2] = data4_s2[2];
	assign data5_s3[0] = data5_s2[0];
	assign data5_s3[1] = data5_s2[1];
	assign data5_s3[2] = data5_s2[2];
	assign data5_s3[3] = data5_s2[3];
	FA F35(.a(data6_s2[0]),.b(data6_s2[1]),.cin(data6_s2[2]),.sum(data6_s3[0]),.cout(data5_s3[4]));
	FA F36(.a(data6_s2[3]),.b(data6_s2[4]),.cin(data6_s2[5]),.sum(data6_s3[1]),.cout(data5_s3[5]));
	FA F37(.a(data7_s2[0]),.b(data7_s2[1]),.cin(data7_s2[2]),.sum(data7_s3[0]),.cout(data6_s3[2]));
	FA F38(.a(data7_s2[3]),.b(data7_s2[4]),.cin(data7_s2[5]),.sum(data7_s3[1]),.cout(data6_s3[3]));
	assign data7_s3[2] = data7_s2[6];
	FA F39(.a(data8_s2[0]),.b(data8_s2[1]),.cin(data8_s2[2]),.sum(data8_s3[0]),.cout(data7_s3[3]));
	assign data8_s3[1] = data8_s2[3];
	HA H4(.a(data9_s2[0]),.cin(data9_s2[1]),.sum(data9_s3[0]),.cout(data8_s3[2]));
	assign data9_s3[1] = data9_s2[2];
	FA F40(.a(data10_s2[0]),.b(data10_s2[1]),.cin(data10_s2[2]),.sum(data10_s3[0]),.cout(data9_s3[2]));
	HA H5(.a(data10_s2[3]),.cin(data10_s2[4]),.sum(data10_s3[1]),.cout(data9_s3[3]));
	FA F41(.a(data11_s2[0]),.b(data11_s2[1]),.cin(data11_s2[2]),.sum(data11_s3[0]),.cout(data10_s3[2]));
	FA F42(.a(data11_s2[3]),.b(data11_s2[4]),.cin(data11_s2[5]),.sum(data11_s3[1]),.cout(data10_s3[3]));
	FA F43(.a(data12_s2[0]),.b(data12_s2[1]),.cin(data12_s2[2]),.sum(data12_s3[0]),.cout(data11_s3[2]));
	FA F44(.a(data12_s2[3]),.b(data12_s2[4]),.cin(data12_s2[5]),.sum(data12_s3[1]),.cout(data11_s3[3]));
	FA F45(.a(data13_s2[0]),.b(data13_s2[1]),.cin(data13_s2[2]),.sum(data13_s3[0]),.cout(data12_s3[2]));
	assign data14_s3[0] = data14_s2[0];
	FA F46(.a(data15_s2[0]),.b(data15_s2[1]),.cin(data15_s2[2]),.sum(data15_s3[0]),.cout(data14_s3[1]));
	assign data15_s3[1] = data15_s2[3];
	assign data15_s3[2] = data15_s2[4];
	assign data16_s3[0] = data16_s2[0];
	assign data17_s3[0] = data17_s2[0];
	assign data18_s3[0] = data18_s2[0];

	//****The 4th stage****
	wire[0:0] data0_s4;
	wire[3:0] data1_s4;
	wire[0:0] data2_s4;
	wire[2:0] data3_s4;
	wire[2:0] data4_s4;
	wire[2:0] data5_s4;
	wire[2:0] data6_s4;
	wire[2:0] data7_s4;
	wire[1:0] data8_s4;
	wire[2:0] data9_s4;
	wire[2:0] data10_s4;
	wire[2:0] data11_s4;
	wire[0:0] data12_s4;
	wire[0:0] data13_s4;
	wire[2:0] data14_s4;
	wire[0:0] data15_s4;
	wire[0:0] data16_s4;
	wire[0:0] data17_s4;
	wire[0:0] data18_s4;
	assign data0_s4[0] = data0_s3[0];
	assign data1_s4[0] = data1_s3[0];
	assign data1_s4[1] = data1_s3[1];
	assign data1_s4[2] = data1_s3[2];
	FA F47(.a(data2_s3[0]),.b(data2_s3[1]),.cin(data2_s3[2]),.sum(data2_s4[0]),.cout(data1_s4[3]));
	assign data3_s4[0] = data3_s3[0];
	assign data3_s4[1] = data3_s3[1];
	FA F48(.a(data4_s3[0]),.b(data4_s3[1]),.cin(data4_s3[2]),.sum(data4_s4[0]),.cout(data3_s4[2]));
	FA F49(.a(data5_s3[0]),.b(data5_s3[1]),.cin(data5_s3[2]),.sum(data5_s4[0]),.cout(data4_s4[1]));
	FA F50(.a(data5_s3[3]),.b(data5_s3[4]),.cin(data5_s3[5]),.sum(data5_s4[1]),.cout(data4_s4[2]));
	FA F51(.a(data6_s3[0]),.b(data6_s3[1]),.cin(data6_s3[2]),.sum(data6_s4[0]),.cout(data5_s4[2]));
	assign data6_s4[1] = data6_s3[3];
	FA F52(.a(data7_s3[0]),.b(data7_s3[1]),.cin(data7_s3[2]),.sum(data7_s4[0]),.cout(data6_s4[2]));
	assign data7_s4[1] = data7_s3[3];
	FA F53(.a(data8_s3[0]),.b(data8_s3[1]),.cin(data8_s3[2]),.sum(data8_s4[0]),.cout(data7_s4[2]));
	FA F54(.a(data9_s3[0]),.b(data9_s3[1]),.cin(data9_s3[2]),.sum(data9_s4[0]),.cout(data8_s4[1]));
	assign data9_s4[1] = data9_s3[3];
	FA F55(.a(data10_s3[0]),.b(data10_s3[1]),.cin(data10_s3[2]),.sum(data10_s4[0]),.cout(data9_s4[2]));
	assign data10_s4[1] = data10_s3[3];
	FA F56(.a(data11_s3[0]),.b(data11_s3[1]),.cin(data11_s3[2]),.sum(data11_s4[0]),.cout(data10_s4[2]));
	assign data11_s4[1] = data11_s3[3];
	FA F57(.a(data12_s3[0]),.b(data12_s3[1]),.cin(data12_s3[2]),.sum(data12_s4[0]),.cout(data11_s4[2]));
	assign data13_s4[0] = data13_s3[0];
	assign data14_s4[0] = data14_s3[0];
	assign data14_s4[1] = data14_s3[1];
	FA F58(.a(data15_s3[0]),.b(data15_s3[1]),.cin(data15_s3[2]),.sum(data15_s4[0]),.cout(data14_s4[2]));
	assign data16_s4[0] = data16_s3[0];
	assign data17_s4[0] = data17_s3[0];
	assign data18_s4[0] = data18_s3[0];

	//****The 5th stage****
	wire[1:0] data0_s5;
	wire[1:0] data1_s5;
	wire[1:0] data2_s5;
	wire[1:0] data3_s5;
	wire[1:0] data4_s5;
	wire[1:0] data5_s5;
	wire[1:0] data6_s5;
	wire[1:0] data7_s5;
	wire[1:0] data8_s5;
	wire[1:0] data9_s5;
	wire[1:0] data10_s5;
	wire[0:0] data11_s5;
	wire[0:0] data12_s5;
	wire[1:0] data13_s5;
	wire[0:0] data14_s5;
	wire[0:0] data15_s5;
	wire[0:0] data16_s5;
	wire[0:0] data17_s5;
	wire[0:0] data18_s5;
	assign data0_s5[0] = data0_s4[0];
	FA F59(.a(data1_s4[0]),.b(data1_s4[1]),.cin(data1_s4[2]),.sum(data1_s5[0]),.cout(data0_s5[1]));
	assign data1_s5[1] = data1_s4[3];
	assign data2_s5[0] = data2_s4[0];
	FA F60(.a(data3_s4[0]),.b(data3_s4[1]),.cin(data3_s4[2]),.sum(data3_s5[0]),.cout(data2_s5[1]));
	FA F61(.a(data4_s4[0]),.b(data4_s4[1]),.cin(data4_s4[2]),.sum(data4_s5[0]),.cout(data3_s5[1]));
	FA F62(.a(data5_s4[0]),.b(data5_s4[1]),.cin(data5_s4[2]),.sum(data5_s5[0]),.cout(data4_s5[1]));
	FA F63(.a(data6_s4[0]),.b(data6_s4[1]),.cin(data6_s4[2]),.sum(data6_s5[0]),.cout(data5_s5[1]));
	FA F64(.a(data7_s4[0]),.b(data7_s4[1]),.cin(data7_s4[2]),.sum(data7_s5[0]),.cout(data6_s5[1]));
	HA H6(.a(data8_s4[0]),.cin(data8_s4[1]),.sum(data8_s5[0]),.cout(data7_s5[1]));
	FA F65(.a(data9_s4[0]),.b(data9_s4[1]),.cin(data9_s4[2]),.sum(data9_s5[0]),.cout(data8_s5[1]));
	FA F66(.a(data10_s4[0]),.b(data10_s4[1]),.cin(data10_s4[2]),.sum(data10_s5[0]),.cout(data9_s5[1]));
	FA F67(.a(data11_s4[0]),.b(data11_s4[1]),.cin(data11_s4[2]),.sum(data11_s5[0]),.cout(data10_s5[1]));
	assign data12_s5[0] = data12_s4[0];
	assign data13_s5[0] = data13_s4[0];
	FA F68(.a(data14_s4[0]),.b(data14_s4[1]),.cin(data14_s4[2]),.sum(data14_s5[0]),.cout(data13_s5[1]));
	assign data15_s5[0] = data15_s4[0];
	assign data16_s5[0] = data16_s4[0];
	assign data17_s5[0] = data17_s4[0];
	assign data18_s5[0] = data18_s4[0];
endmodule
